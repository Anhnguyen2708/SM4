library verilog;
use verilog.vl_types.all;
entity sm4_top_vlg_vec_tst is
end sm4_top_vlg_vec_tst;
